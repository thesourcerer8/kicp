VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Matrix_Multiplication
  CLASS BLOCK ;
  FOREIGN Matrix_Multiplication ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1760.000 ;
  PIN addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END addr_o[0]
  PIN addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.910 0.000 1020.190 4.000 ;
    END
  END addr_o[10]
  PIN addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.330 0.000 1101.610 4.000 ;
    END
  END addr_o[11]
  PIN addr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.750 0.000 1183.030 4.000 ;
    END
  END addr_o[12]
  PIN addr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.170 0.000 1264.450 4.000 ;
    END
  END addr_o[13]
  PIN addr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.590 0.000 1345.870 4.000 ;
    END
  END addr_o[14]
  PIN addr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.010 0.000 1427.290 4.000 ;
    END
  END addr_o[15]
  PIN addr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.430 0.000 1508.710 4.000 ;
    END
  END addr_o[16]
  PIN addr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.850 0.000 1590.130 4.000 ;
    END
  END addr_o[17]
  PIN addr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.270 0.000 1671.550 4.000 ;
    END
  END addr_o[18]
  PIN addr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.690 0.000 1752.970 4.000 ;
    END
  END addr_o[19]
  PIN addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END addr_o[1]
  PIN addr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.110 0.000 1834.390 4.000 ;
    END
  END addr_o[20]
  PIN addr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.530 0.000 1915.810 4.000 ;
    END
  END addr_o[21]
  PIN addr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1996.950 0.000 1997.230 4.000 ;
    END
  END addr_o[22]
  PIN addr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2078.370 0.000 2078.650 4.000 ;
    END
  END addr_o[23]
  PIN addr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2159.790 0.000 2160.070 4.000 ;
    END
  END addr_o[24]
  PIN addr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2241.210 0.000 2241.490 4.000 ;
    END
  END addr_o[25]
  PIN addr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2322.630 0.000 2322.910 4.000 ;
    END
  END addr_o[26]
  PIN addr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2404.050 0.000 2404.330 4.000 ;
    END
  END addr_o[27]
  PIN addr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.470 0.000 2485.750 4.000 ;
    END
  END addr_o[28]
  PIN addr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2566.890 0.000 2567.170 4.000 ;
    END
  END addr_o[29]
  PIN addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END addr_o[2]
  PIN addr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2648.310 0.000 2648.590 4.000 ;
    END
  END addr_o[30]
  PIN addr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2729.730 0.000 2730.010 4.000 ;
    END
  END addr_o[31]
  PIN addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END addr_o[3]
  PIN addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END addr_o[4]
  PIN addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 0.000 613.090 4.000 ;
    END
  END addr_o[5]
  PIN addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END addr_o[6]
  PIN addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 0.000 775.930 4.000 ;
    END
  END addr_o[7]
  PIN addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.070 0.000 857.350 4.000 ;
    END
  END addr_o[8]
  PIN addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.490 0.000 938.770 4.000 ;
    END
  END addr_o[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END clk
  PIN data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END data_i[0]
  PIN data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.050 0.000 1047.330 4.000 ;
    END
  END data_i[10]
  PIN data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.470 0.000 1128.750 4.000 ;
    END
  END data_i[11]
  PIN data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.890 0.000 1210.170 4.000 ;
    END
  END data_i[12]
  PIN data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 0.000 1291.590 4.000 ;
    END
  END data_i[13]
  PIN data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1372.730 0.000 1373.010 4.000 ;
    END
  END data_i[14]
  PIN data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.150 0.000 1454.430 4.000 ;
    END
  END data_i[15]
  PIN data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.570 0.000 1535.850 4.000 ;
    END
  END data_i[16]
  PIN data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.990 0.000 1617.270 4.000 ;
    END
  END data_i[17]
  PIN data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1698.410 0.000 1698.690 4.000 ;
    END
  END data_i[18]
  PIN data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1779.830 0.000 1780.110 4.000 ;
    END
  END data_i[19]
  PIN data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END data_i[1]
  PIN data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.250 0.000 1861.530 4.000 ;
    END
  END data_i[20]
  PIN data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1942.670 0.000 1942.950 4.000 ;
    END
  END data_i[21]
  PIN data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2024.090 0.000 2024.370 4.000 ;
    END
  END data_i[22]
  PIN data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2105.510 0.000 2105.790 4.000 ;
    END
  END data_i[23]
  PIN data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2186.930 0.000 2187.210 4.000 ;
    END
  END data_i[24]
  PIN data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2268.350 0.000 2268.630 4.000 ;
    END
  END data_i[25]
  PIN data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2349.770 0.000 2350.050 4.000 ;
    END
  END data_i[26]
  PIN data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.190 0.000 2431.470 4.000 ;
    END
  END data_i[27]
  PIN data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2512.610 0.000 2512.890 4.000 ;
    END
  END data_i[28]
  PIN data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2594.030 0.000 2594.310 4.000 ;
    END
  END data_i[29]
  PIN data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END data_i[2]
  PIN data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2675.450 0.000 2675.730 4.000 ;
    END
  END data_i[30]
  PIN data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2756.870 0.000 2757.150 4.000 ;
    END
  END data_i[31]
  PIN data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 0.000 477.390 4.000 ;
    END
  END data_i[3]
  PIN data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 0.000 558.810 4.000 ;
    END
  END data_i[4]
  PIN data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 0.000 640.230 4.000 ;
    END
  END data_i[5]
  PIN data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 0.000 721.650 4.000 ;
    END
  END data_i[6]
  PIN data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.790 0.000 803.070 4.000 ;
    END
  END data_i[7]
  PIN data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.210 0.000 884.490 4.000 ;
    END
  END data_i[8]
  PIN data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.630 0.000 965.910 4.000 ;
    END
  END data_i[9]
  PIN data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END data_o[0]
  PIN data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1074.190 0.000 1074.470 4.000 ;
    END
  END data_o[10]
  PIN data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.610 0.000 1155.890 4.000 ;
    END
  END data_o[11]
  PIN data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.030 0.000 1237.310 4.000 ;
    END
  END data_o[12]
  PIN data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.450 0.000 1318.730 4.000 ;
    END
  END data_o[13]
  PIN data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.870 0.000 1400.150 4.000 ;
    END
  END data_o[14]
  PIN data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.290 0.000 1481.570 4.000 ;
    END
  END data_o[15]
  PIN data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1562.710 0.000 1562.990 4.000 ;
    END
  END data_o[16]
  PIN data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1644.130 0.000 1644.410 4.000 ;
    END
  END data_o[17]
  PIN data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1725.550 0.000 1725.830 4.000 ;
    END
  END data_o[18]
  PIN data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1806.970 0.000 1807.250 4.000 ;
    END
  END data_o[19]
  PIN data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END data_o[1]
  PIN data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.390 0.000 1888.670 4.000 ;
    END
  END data_o[20]
  PIN data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1969.810 0.000 1970.090 4.000 ;
    END
  END data_o[21]
  PIN data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2051.230 0.000 2051.510 4.000 ;
    END
  END data_o[22]
  PIN data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2132.650 0.000 2132.930 4.000 ;
    END
  END data_o[23]
  PIN data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2214.070 0.000 2214.350 4.000 ;
    END
  END data_o[24]
  PIN data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.490 0.000 2295.770 4.000 ;
    END
  END data_o[25]
  PIN data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2376.910 0.000 2377.190 4.000 ;
    END
  END data_o[26]
  PIN data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2458.330 0.000 2458.610 4.000 ;
    END
  END data_o[27]
  PIN data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2539.750 0.000 2540.030 4.000 ;
    END
  END data_o[28]
  PIN data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.170 0.000 2621.450 4.000 ;
    END
  END data_o[29]
  PIN data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 4.000 ;
    END
  END data_o[2]
  PIN data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2702.590 0.000 2702.870 4.000 ;
    END
  END data_o[30]
  PIN data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2784.010 0.000 2784.290 4.000 ;
    END
  END data_o[31]
  PIN data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 0.000 504.530 4.000 ;
    END
  END data_o[3]
  PIN data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 0.000 585.950 4.000 ;
    END
  END data_o[4]
  PIN data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END data_o[5]
  PIN data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.510 0.000 748.790 4.000 ;
    END
  END data_o[6]
  PIN data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.930 0.000 830.210 4.000 ;
    END
  END data_o[7]
  PIN data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 0.000 911.630 4.000 ;
    END
  END data_o[8]
  PIN data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.770 0.000 993.050 4.000 ;
    END
  END data_o[9]
  PIN done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END done
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END enable
  PIN mem_opdone
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END mem_opdone
  PIN mem_operation[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END mem_operation[0]
  PIN mem_operation[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END mem_operation[1]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2785.840 10.640 2787.440 1749.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 1749.200 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 1747.545 2794.230 1749.150 ;
        RECT 5.330 1742.105 2794.230 1744.935 ;
        RECT 5.330 1736.665 2794.230 1739.495 ;
        RECT 5.330 1731.225 2794.230 1734.055 ;
        RECT 5.330 1725.785 2794.230 1728.615 ;
        RECT 5.330 1720.345 2794.230 1723.175 ;
        RECT 5.330 1714.905 2794.230 1717.735 ;
        RECT 5.330 1709.465 2794.230 1712.295 ;
        RECT 5.330 1704.025 2794.230 1706.855 ;
        RECT 5.330 1698.585 2794.230 1701.415 ;
        RECT 5.330 1693.145 2794.230 1695.975 ;
        RECT 5.330 1687.705 2794.230 1690.535 ;
        RECT 5.330 1682.265 2794.230 1685.095 ;
        RECT 5.330 1676.825 2794.230 1679.655 ;
        RECT 5.330 1671.385 2794.230 1674.215 ;
        RECT 5.330 1665.945 2794.230 1668.775 ;
        RECT 5.330 1660.505 2794.230 1663.335 ;
        RECT 5.330 1655.065 2794.230 1657.895 ;
        RECT 5.330 1649.625 2794.230 1652.455 ;
        RECT 5.330 1644.185 2794.230 1647.015 ;
        RECT 5.330 1638.745 2794.230 1641.575 ;
        RECT 5.330 1633.305 2794.230 1636.135 ;
        RECT 5.330 1627.865 2794.230 1630.695 ;
        RECT 5.330 1622.425 2794.230 1625.255 ;
        RECT 5.330 1616.985 2794.230 1619.815 ;
        RECT 5.330 1611.545 2794.230 1614.375 ;
        RECT 5.330 1606.105 2794.230 1608.935 ;
        RECT 5.330 1600.665 2794.230 1603.495 ;
        RECT 5.330 1595.225 2794.230 1598.055 ;
        RECT 5.330 1589.785 2794.230 1592.615 ;
        RECT 5.330 1584.345 2794.230 1587.175 ;
        RECT 5.330 1578.905 2794.230 1581.735 ;
        RECT 5.330 1573.465 2794.230 1576.295 ;
        RECT 5.330 1568.025 2794.230 1570.855 ;
        RECT 5.330 1562.585 2794.230 1565.415 ;
        RECT 5.330 1557.145 2794.230 1559.975 ;
        RECT 5.330 1551.705 2794.230 1554.535 ;
        RECT 5.330 1546.265 2794.230 1549.095 ;
        RECT 5.330 1540.825 2794.230 1543.655 ;
        RECT 5.330 1535.385 2794.230 1538.215 ;
        RECT 5.330 1529.945 2794.230 1532.775 ;
        RECT 5.330 1524.505 2794.230 1527.335 ;
        RECT 5.330 1519.065 2794.230 1521.895 ;
        RECT 5.330 1513.625 2794.230 1516.455 ;
        RECT 5.330 1508.185 2794.230 1511.015 ;
        RECT 5.330 1502.745 2794.230 1505.575 ;
        RECT 5.330 1497.305 2794.230 1500.135 ;
        RECT 5.330 1491.865 2794.230 1494.695 ;
        RECT 5.330 1486.425 2794.230 1489.255 ;
        RECT 5.330 1480.985 2794.230 1483.815 ;
        RECT 5.330 1475.545 2794.230 1478.375 ;
        RECT 5.330 1470.105 2794.230 1472.935 ;
        RECT 5.330 1464.665 2794.230 1467.495 ;
        RECT 5.330 1459.225 2794.230 1462.055 ;
        RECT 5.330 1453.785 2794.230 1456.615 ;
        RECT 5.330 1448.345 2794.230 1451.175 ;
        RECT 5.330 1442.905 2794.230 1445.735 ;
        RECT 5.330 1437.465 2794.230 1440.295 ;
        RECT 5.330 1432.025 2794.230 1434.855 ;
        RECT 5.330 1426.585 2794.230 1429.415 ;
        RECT 5.330 1421.145 2794.230 1423.975 ;
        RECT 5.330 1415.705 2794.230 1418.535 ;
        RECT 5.330 1410.265 2794.230 1413.095 ;
        RECT 5.330 1404.825 2794.230 1407.655 ;
        RECT 5.330 1399.385 2794.230 1402.215 ;
        RECT 5.330 1393.945 2794.230 1396.775 ;
        RECT 5.330 1388.505 2794.230 1391.335 ;
        RECT 5.330 1383.065 2794.230 1385.895 ;
        RECT 5.330 1377.625 2794.230 1380.455 ;
        RECT 5.330 1372.185 2794.230 1375.015 ;
        RECT 5.330 1366.745 2794.230 1369.575 ;
        RECT 5.330 1361.305 2794.230 1364.135 ;
        RECT 5.330 1355.865 2794.230 1358.695 ;
        RECT 5.330 1350.425 2794.230 1353.255 ;
        RECT 5.330 1344.985 2794.230 1347.815 ;
        RECT 5.330 1339.545 2794.230 1342.375 ;
        RECT 5.330 1334.105 2794.230 1336.935 ;
        RECT 5.330 1328.665 2794.230 1331.495 ;
        RECT 5.330 1323.225 2794.230 1326.055 ;
        RECT 5.330 1317.785 2794.230 1320.615 ;
        RECT 5.330 1312.345 2794.230 1315.175 ;
        RECT 5.330 1306.905 2794.230 1309.735 ;
        RECT 5.330 1301.465 2794.230 1304.295 ;
        RECT 5.330 1296.025 2794.230 1298.855 ;
        RECT 5.330 1290.585 2794.230 1293.415 ;
        RECT 5.330 1285.145 2794.230 1287.975 ;
        RECT 5.330 1279.705 2794.230 1282.535 ;
        RECT 5.330 1274.265 2794.230 1277.095 ;
        RECT 5.330 1268.825 2794.230 1271.655 ;
        RECT 5.330 1263.385 2794.230 1266.215 ;
        RECT 5.330 1257.945 2794.230 1260.775 ;
        RECT 5.330 1252.505 2794.230 1255.335 ;
        RECT 5.330 1247.065 2794.230 1249.895 ;
        RECT 5.330 1241.625 2794.230 1244.455 ;
        RECT 5.330 1236.185 2794.230 1239.015 ;
        RECT 5.330 1230.745 2794.230 1233.575 ;
        RECT 5.330 1225.305 2794.230 1228.135 ;
        RECT 5.330 1219.865 2794.230 1222.695 ;
        RECT 5.330 1214.425 2794.230 1217.255 ;
        RECT 5.330 1208.985 2794.230 1211.815 ;
        RECT 5.330 1203.545 2794.230 1206.375 ;
        RECT 5.330 1198.105 2794.230 1200.935 ;
        RECT 5.330 1192.665 2794.230 1195.495 ;
        RECT 5.330 1187.225 2794.230 1190.055 ;
        RECT 5.330 1181.785 2794.230 1184.615 ;
        RECT 5.330 1176.345 2794.230 1179.175 ;
        RECT 5.330 1170.905 2794.230 1173.735 ;
        RECT 5.330 1165.465 2794.230 1168.295 ;
        RECT 5.330 1160.025 2794.230 1162.855 ;
        RECT 5.330 1154.585 2794.230 1157.415 ;
        RECT 5.330 1149.145 2794.230 1151.975 ;
        RECT 5.330 1143.705 2794.230 1146.535 ;
        RECT 5.330 1138.265 2794.230 1141.095 ;
        RECT 5.330 1132.825 2794.230 1135.655 ;
        RECT 5.330 1127.385 2794.230 1130.215 ;
        RECT 5.330 1121.945 2794.230 1124.775 ;
        RECT 5.330 1116.505 2794.230 1119.335 ;
        RECT 5.330 1111.065 2794.230 1113.895 ;
        RECT 5.330 1105.625 2794.230 1108.455 ;
        RECT 5.330 1100.185 2794.230 1103.015 ;
        RECT 5.330 1094.745 2794.230 1097.575 ;
        RECT 5.330 1089.305 2794.230 1092.135 ;
        RECT 5.330 1083.865 2794.230 1086.695 ;
        RECT 5.330 1078.425 2794.230 1081.255 ;
        RECT 5.330 1072.985 2794.230 1075.815 ;
        RECT 5.330 1067.545 2794.230 1070.375 ;
        RECT 5.330 1062.105 2794.230 1064.935 ;
        RECT 5.330 1056.665 2794.230 1059.495 ;
        RECT 5.330 1051.225 2794.230 1054.055 ;
        RECT 5.330 1045.785 2794.230 1048.615 ;
        RECT 5.330 1040.345 2794.230 1043.175 ;
        RECT 5.330 1034.905 2794.230 1037.735 ;
        RECT 5.330 1029.465 2794.230 1032.295 ;
        RECT 5.330 1024.025 2794.230 1026.855 ;
        RECT 5.330 1018.585 2794.230 1021.415 ;
        RECT 5.330 1013.145 2794.230 1015.975 ;
        RECT 5.330 1007.705 2794.230 1010.535 ;
        RECT 5.330 1002.265 2794.230 1005.095 ;
        RECT 5.330 996.825 2794.230 999.655 ;
        RECT 5.330 991.385 2794.230 994.215 ;
        RECT 5.330 985.945 2794.230 988.775 ;
        RECT 5.330 980.505 2794.230 983.335 ;
        RECT 5.330 975.065 2794.230 977.895 ;
        RECT 5.330 969.625 2794.230 972.455 ;
        RECT 5.330 964.185 2794.230 967.015 ;
        RECT 5.330 958.745 2794.230 961.575 ;
        RECT 5.330 953.305 2794.230 956.135 ;
        RECT 5.330 947.865 2794.230 950.695 ;
        RECT 5.330 942.425 2794.230 945.255 ;
        RECT 5.330 936.985 2794.230 939.815 ;
        RECT 5.330 931.545 2794.230 934.375 ;
        RECT 5.330 926.105 2794.230 928.935 ;
        RECT 5.330 920.665 2794.230 923.495 ;
        RECT 5.330 915.225 2794.230 918.055 ;
        RECT 5.330 909.785 2794.230 912.615 ;
        RECT 5.330 904.345 2794.230 907.175 ;
        RECT 5.330 898.905 2794.230 901.735 ;
        RECT 5.330 893.465 2794.230 896.295 ;
        RECT 5.330 888.025 2794.230 890.855 ;
        RECT 5.330 882.585 2794.230 885.415 ;
        RECT 5.330 877.145 2794.230 879.975 ;
        RECT 5.330 871.705 2794.230 874.535 ;
        RECT 5.330 866.265 2794.230 869.095 ;
        RECT 5.330 860.825 2794.230 863.655 ;
        RECT 5.330 855.385 2794.230 858.215 ;
        RECT 5.330 849.945 2794.230 852.775 ;
        RECT 5.330 844.505 2794.230 847.335 ;
        RECT 5.330 839.065 2794.230 841.895 ;
        RECT 5.330 833.625 2794.230 836.455 ;
        RECT 5.330 828.185 2794.230 831.015 ;
        RECT 5.330 822.745 2794.230 825.575 ;
        RECT 5.330 817.305 2794.230 820.135 ;
        RECT 5.330 811.865 2794.230 814.695 ;
        RECT 5.330 806.425 2794.230 809.255 ;
        RECT 5.330 800.985 2794.230 803.815 ;
        RECT 5.330 795.545 2794.230 798.375 ;
        RECT 5.330 790.105 2794.230 792.935 ;
        RECT 5.330 784.665 2794.230 787.495 ;
        RECT 5.330 779.225 2794.230 782.055 ;
        RECT 5.330 773.785 2794.230 776.615 ;
        RECT 5.330 768.345 2794.230 771.175 ;
        RECT 5.330 762.905 2794.230 765.735 ;
        RECT 5.330 757.465 2794.230 760.295 ;
        RECT 5.330 752.025 2794.230 754.855 ;
        RECT 5.330 746.585 2794.230 749.415 ;
        RECT 5.330 741.145 2794.230 743.975 ;
        RECT 5.330 735.705 2794.230 738.535 ;
        RECT 5.330 730.265 2794.230 733.095 ;
        RECT 5.330 724.825 2794.230 727.655 ;
        RECT 5.330 719.385 2794.230 722.215 ;
        RECT 5.330 713.945 2794.230 716.775 ;
        RECT 5.330 708.505 2794.230 711.335 ;
        RECT 5.330 703.065 2794.230 705.895 ;
        RECT 5.330 697.625 2794.230 700.455 ;
        RECT 5.330 692.185 2794.230 695.015 ;
        RECT 5.330 686.745 2794.230 689.575 ;
        RECT 5.330 681.305 2794.230 684.135 ;
        RECT 5.330 675.865 2794.230 678.695 ;
        RECT 5.330 670.425 2794.230 673.255 ;
        RECT 5.330 664.985 2794.230 667.815 ;
        RECT 5.330 659.545 2794.230 662.375 ;
        RECT 5.330 654.105 2794.230 656.935 ;
        RECT 5.330 648.665 2794.230 651.495 ;
        RECT 5.330 643.225 2794.230 646.055 ;
        RECT 5.330 637.785 2794.230 640.615 ;
        RECT 5.330 632.345 2794.230 635.175 ;
        RECT 5.330 626.905 2794.230 629.735 ;
        RECT 5.330 621.465 2794.230 624.295 ;
        RECT 5.330 616.025 2794.230 618.855 ;
        RECT 5.330 610.585 2794.230 613.415 ;
        RECT 5.330 605.145 2794.230 607.975 ;
        RECT 5.330 599.705 2794.230 602.535 ;
        RECT 5.330 594.265 2794.230 597.095 ;
        RECT 5.330 588.825 2794.230 591.655 ;
        RECT 5.330 583.385 2794.230 586.215 ;
        RECT 5.330 577.945 2794.230 580.775 ;
        RECT 5.330 572.505 2794.230 575.335 ;
        RECT 5.330 567.065 2794.230 569.895 ;
        RECT 5.330 561.625 2794.230 564.455 ;
        RECT 5.330 556.185 2794.230 559.015 ;
        RECT 5.330 550.745 2794.230 553.575 ;
        RECT 5.330 545.305 2794.230 548.135 ;
        RECT 5.330 539.865 2794.230 542.695 ;
        RECT 5.330 534.425 2794.230 537.255 ;
        RECT 5.330 528.985 2794.230 531.815 ;
        RECT 5.330 523.545 2794.230 526.375 ;
        RECT 5.330 518.105 2794.230 520.935 ;
        RECT 5.330 512.665 2794.230 515.495 ;
        RECT 5.330 507.225 2794.230 510.055 ;
        RECT 5.330 501.785 2794.230 504.615 ;
        RECT 5.330 496.345 2794.230 499.175 ;
        RECT 5.330 490.905 2794.230 493.735 ;
        RECT 5.330 485.465 2794.230 488.295 ;
        RECT 5.330 480.025 2794.230 482.855 ;
        RECT 5.330 474.585 2794.230 477.415 ;
        RECT 5.330 469.145 2794.230 471.975 ;
        RECT 5.330 463.705 2794.230 466.535 ;
        RECT 5.330 458.265 2794.230 461.095 ;
        RECT 5.330 452.825 2794.230 455.655 ;
        RECT 5.330 447.385 2794.230 450.215 ;
        RECT 5.330 441.945 2794.230 444.775 ;
        RECT 5.330 436.505 2794.230 439.335 ;
        RECT 5.330 431.065 2794.230 433.895 ;
        RECT 5.330 425.625 2794.230 428.455 ;
        RECT 5.330 420.185 2794.230 423.015 ;
        RECT 5.330 414.745 2794.230 417.575 ;
        RECT 5.330 409.305 2794.230 412.135 ;
        RECT 5.330 403.865 2794.230 406.695 ;
        RECT 5.330 398.425 2794.230 401.255 ;
        RECT 5.330 392.985 2794.230 395.815 ;
        RECT 5.330 387.545 2794.230 390.375 ;
        RECT 5.330 382.105 2794.230 384.935 ;
        RECT 5.330 376.665 2794.230 379.495 ;
        RECT 5.330 371.225 2794.230 374.055 ;
        RECT 5.330 365.785 2794.230 368.615 ;
        RECT 5.330 360.345 2794.230 363.175 ;
        RECT 5.330 354.905 2794.230 357.735 ;
        RECT 5.330 349.465 2794.230 352.295 ;
        RECT 5.330 344.025 2794.230 346.855 ;
        RECT 5.330 338.585 2794.230 341.415 ;
        RECT 5.330 333.145 2794.230 335.975 ;
        RECT 5.330 327.705 2794.230 330.535 ;
        RECT 5.330 322.265 2794.230 325.095 ;
        RECT 5.330 316.825 2794.230 319.655 ;
        RECT 5.330 311.385 2794.230 314.215 ;
        RECT 5.330 305.945 2794.230 308.775 ;
        RECT 5.330 300.505 2794.230 303.335 ;
        RECT 5.330 295.065 2794.230 297.895 ;
        RECT 5.330 289.625 2794.230 292.455 ;
        RECT 5.330 284.185 2794.230 287.015 ;
        RECT 5.330 278.745 2794.230 281.575 ;
        RECT 5.330 273.305 2794.230 276.135 ;
        RECT 5.330 267.865 2794.230 270.695 ;
        RECT 5.330 262.425 2794.230 265.255 ;
        RECT 5.330 256.985 2794.230 259.815 ;
        RECT 5.330 251.545 2794.230 254.375 ;
        RECT 5.330 246.105 2794.230 248.935 ;
        RECT 5.330 240.665 2794.230 243.495 ;
        RECT 5.330 235.225 2794.230 238.055 ;
        RECT 5.330 229.785 2794.230 232.615 ;
        RECT 5.330 224.345 2794.230 227.175 ;
        RECT 5.330 218.905 2794.230 221.735 ;
        RECT 5.330 213.465 2794.230 216.295 ;
        RECT 5.330 208.025 2794.230 210.855 ;
        RECT 5.330 202.585 2794.230 205.415 ;
        RECT 5.330 197.145 2794.230 199.975 ;
        RECT 5.330 191.705 2794.230 194.535 ;
        RECT 5.330 186.265 2794.230 189.095 ;
        RECT 5.330 180.825 2794.230 183.655 ;
        RECT 5.330 175.385 2794.230 178.215 ;
        RECT 5.330 169.945 2794.230 172.775 ;
        RECT 5.330 164.505 2794.230 167.335 ;
        RECT 5.330 159.065 2794.230 161.895 ;
        RECT 5.330 153.625 2794.230 156.455 ;
        RECT 5.330 148.185 2794.230 151.015 ;
        RECT 5.330 142.745 2794.230 145.575 ;
        RECT 5.330 137.305 2794.230 140.135 ;
        RECT 5.330 131.865 2794.230 134.695 ;
        RECT 5.330 126.425 2794.230 129.255 ;
        RECT 5.330 120.985 2794.230 123.815 ;
        RECT 5.330 115.545 2794.230 118.375 ;
        RECT 5.330 110.105 2794.230 112.935 ;
        RECT 5.330 104.665 2794.230 107.495 ;
        RECT 5.330 99.225 2794.230 102.055 ;
        RECT 5.330 93.785 2794.230 96.615 ;
        RECT 5.330 88.345 2794.230 91.175 ;
        RECT 5.330 82.905 2794.230 85.735 ;
        RECT 5.330 77.465 2794.230 80.295 ;
        RECT 5.330 72.025 2794.230 74.855 ;
        RECT 5.330 66.585 2794.230 69.415 ;
        RECT 5.330 61.145 2794.230 63.975 ;
        RECT 5.330 55.705 2794.230 58.535 ;
        RECT 5.330 50.265 2794.230 53.095 ;
        RECT 5.330 44.825 2794.230 47.655 ;
        RECT 5.330 39.385 2794.230 42.215 ;
        RECT 5.330 33.945 2794.230 36.775 ;
        RECT 5.330 28.505 2794.230 31.335 ;
        RECT 5.330 23.065 2794.230 25.895 ;
        RECT 5.330 17.625 2794.230 20.455 ;
        RECT 5.330 12.185 2794.230 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 2794.040 1749.045 ;
      LAYER met1 ;
        RECT 5.520 0.380 2794.040 1749.200 ;
      LAYER met2 ;
        RECT 21.070 4.280 2787.410 1749.145 ;
        RECT 21.070 0.350 42.590 4.280 ;
        RECT 43.430 0.350 69.730 4.280 ;
        RECT 70.570 0.350 96.870 4.280 ;
        RECT 97.710 0.350 124.010 4.280 ;
        RECT 124.850 0.350 151.150 4.280 ;
        RECT 151.990 0.350 178.290 4.280 ;
        RECT 179.130 0.350 205.430 4.280 ;
        RECT 206.270 0.350 232.570 4.280 ;
        RECT 233.410 0.350 259.710 4.280 ;
        RECT 260.550 0.350 286.850 4.280 ;
        RECT 287.690 0.350 313.990 4.280 ;
        RECT 314.830 0.350 341.130 4.280 ;
        RECT 341.970 0.350 368.270 4.280 ;
        RECT 369.110 0.350 395.410 4.280 ;
        RECT 396.250 0.350 422.550 4.280 ;
        RECT 423.390 0.350 449.690 4.280 ;
        RECT 450.530 0.350 476.830 4.280 ;
        RECT 477.670 0.350 503.970 4.280 ;
        RECT 504.810 0.350 531.110 4.280 ;
        RECT 531.950 0.350 558.250 4.280 ;
        RECT 559.090 0.350 585.390 4.280 ;
        RECT 586.230 0.350 612.530 4.280 ;
        RECT 613.370 0.350 639.670 4.280 ;
        RECT 640.510 0.350 666.810 4.280 ;
        RECT 667.650 0.350 693.950 4.280 ;
        RECT 694.790 0.350 721.090 4.280 ;
        RECT 721.930 0.350 748.230 4.280 ;
        RECT 749.070 0.350 775.370 4.280 ;
        RECT 776.210 0.350 802.510 4.280 ;
        RECT 803.350 0.350 829.650 4.280 ;
        RECT 830.490 0.350 856.790 4.280 ;
        RECT 857.630 0.350 883.930 4.280 ;
        RECT 884.770 0.350 911.070 4.280 ;
        RECT 911.910 0.350 938.210 4.280 ;
        RECT 939.050 0.350 965.350 4.280 ;
        RECT 966.190 0.350 992.490 4.280 ;
        RECT 993.330 0.350 1019.630 4.280 ;
        RECT 1020.470 0.350 1046.770 4.280 ;
        RECT 1047.610 0.350 1073.910 4.280 ;
        RECT 1074.750 0.350 1101.050 4.280 ;
        RECT 1101.890 0.350 1128.190 4.280 ;
        RECT 1129.030 0.350 1155.330 4.280 ;
        RECT 1156.170 0.350 1182.470 4.280 ;
        RECT 1183.310 0.350 1209.610 4.280 ;
        RECT 1210.450 0.350 1236.750 4.280 ;
        RECT 1237.590 0.350 1263.890 4.280 ;
        RECT 1264.730 0.350 1291.030 4.280 ;
        RECT 1291.870 0.350 1318.170 4.280 ;
        RECT 1319.010 0.350 1345.310 4.280 ;
        RECT 1346.150 0.350 1372.450 4.280 ;
        RECT 1373.290 0.350 1399.590 4.280 ;
        RECT 1400.430 0.350 1426.730 4.280 ;
        RECT 1427.570 0.350 1453.870 4.280 ;
        RECT 1454.710 0.350 1481.010 4.280 ;
        RECT 1481.850 0.350 1508.150 4.280 ;
        RECT 1508.990 0.350 1535.290 4.280 ;
        RECT 1536.130 0.350 1562.430 4.280 ;
        RECT 1563.270 0.350 1589.570 4.280 ;
        RECT 1590.410 0.350 1616.710 4.280 ;
        RECT 1617.550 0.350 1643.850 4.280 ;
        RECT 1644.690 0.350 1670.990 4.280 ;
        RECT 1671.830 0.350 1698.130 4.280 ;
        RECT 1698.970 0.350 1725.270 4.280 ;
        RECT 1726.110 0.350 1752.410 4.280 ;
        RECT 1753.250 0.350 1779.550 4.280 ;
        RECT 1780.390 0.350 1806.690 4.280 ;
        RECT 1807.530 0.350 1833.830 4.280 ;
        RECT 1834.670 0.350 1860.970 4.280 ;
        RECT 1861.810 0.350 1888.110 4.280 ;
        RECT 1888.950 0.350 1915.250 4.280 ;
        RECT 1916.090 0.350 1942.390 4.280 ;
        RECT 1943.230 0.350 1969.530 4.280 ;
        RECT 1970.370 0.350 1996.670 4.280 ;
        RECT 1997.510 0.350 2023.810 4.280 ;
        RECT 2024.650 0.350 2050.950 4.280 ;
        RECT 2051.790 0.350 2078.090 4.280 ;
        RECT 2078.930 0.350 2105.230 4.280 ;
        RECT 2106.070 0.350 2132.370 4.280 ;
        RECT 2133.210 0.350 2159.510 4.280 ;
        RECT 2160.350 0.350 2186.650 4.280 ;
        RECT 2187.490 0.350 2213.790 4.280 ;
        RECT 2214.630 0.350 2240.930 4.280 ;
        RECT 2241.770 0.350 2268.070 4.280 ;
        RECT 2268.910 0.350 2295.210 4.280 ;
        RECT 2296.050 0.350 2322.350 4.280 ;
        RECT 2323.190 0.350 2349.490 4.280 ;
        RECT 2350.330 0.350 2376.630 4.280 ;
        RECT 2377.470 0.350 2403.770 4.280 ;
        RECT 2404.610 0.350 2430.910 4.280 ;
        RECT 2431.750 0.350 2458.050 4.280 ;
        RECT 2458.890 0.350 2485.190 4.280 ;
        RECT 2486.030 0.350 2512.330 4.280 ;
        RECT 2513.170 0.350 2539.470 4.280 ;
        RECT 2540.310 0.350 2566.610 4.280 ;
        RECT 2567.450 0.350 2593.750 4.280 ;
        RECT 2594.590 0.350 2620.890 4.280 ;
        RECT 2621.730 0.350 2648.030 4.280 ;
        RECT 2648.870 0.350 2675.170 4.280 ;
        RECT 2676.010 0.350 2702.310 4.280 ;
        RECT 2703.150 0.350 2729.450 4.280 ;
        RECT 2730.290 0.350 2756.590 4.280 ;
        RECT 2757.430 0.350 2783.730 4.280 ;
        RECT 2784.570 0.350 2787.410 4.280 ;
      LAYER met3 ;
        RECT 21.050 10.715 2787.430 1749.125 ;
  END
END Matrix_Multiplication
END LIBRARY

