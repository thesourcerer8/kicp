magic
tech sky130A
magscale 1 2
timestamp 1685803793
<< nwell >>
rect 1066 349509 558846 349830
rect 1066 348421 558846 348987
rect 1066 347333 558846 347899
rect 1066 346245 558846 346811
rect 1066 345157 558846 345723
rect 1066 344069 558846 344635
rect 1066 342981 558846 343547
rect 1066 341893 558846 342459
rect 1066 340805 558846 341371
rect 1066 339717 558846 340283
rect 1066 338629 558846 339195
rect 1066 337541 558846 338107
rect 1066 336453 558846 337019
rect 1066 335365 558846 335931
rect 1066 334277 558846 334843
rect 1066 333189 558846 333755
rect 1066 332101 558846 332667
rect 1066 331013 558846 331579
rect 1066 329925 558846 330491
rect 1066 328837 558846 329403
rect 1066 327749 558846 328315
rect 1066 326661 558846 327227
rect 1066 325573 558846 326139
rect 1066 324485 558846 325051
rect 1066 323397 558846 323963
rect 1066 322309 558846 322875
rect 1066 321221 558846 321787
rect 1066 320133 558846 320699
rect 1066 319045 558846 319611
rect 1066 317957 558846 318523
rect 1066 316869 558846 317435
rect 1066 315781 558846 316347
rect 1066 314693 558846 315259
rect 1066 313605 558846 314171
rect 1066 312517 558846 313083
rect 1066 311429 558846 311995
rect 1066 310341 558846 310907
rect 1066 309253 558846 309819
rect 1066 308165 558846 308731
rect 1066 307077 558846 307643
rect 1066 305989 558846 306555
rect 1066 304901 558846 305467
rect 1066 303813 558846 304379
rect 1066 302725 558846 303291
rect 1066 301637 558846 302203
rect 1066 300549 558846 301115
rect 1066 299461 558846 300027
rect 1066 298373 558846 298939
rect 1066 297285 558846 297851
rect 1066 296197 558846 296763
rect 1066 295109 558846 295675
rect 1066 294021 558846 294587
rect 1066 292933 558846 293499
rect 1066 291845 558846 292411
rect 1066 290757 558846 291323
rect 1066 289669 558846 290235
rect 1066 288581 558846 289147
rect 1066 287493 558846 288059
rect 1066 286405 558846 286971
rect 1066 285317 558846 285883
rect 1066 284229 558846 284795
rect 1066 283141 558846 283707
rect 1066 282053 558846 282619
rect 1066 280965 558846 281531
rect 1066 279877 558846 280443
rect 1066 278789 558846 279355
rect 1066 277701 558846 278267
rect 1066 276613 558846 277179
rect 1066 275525 558846 276091
rect 1066 274437 558846 275003
rect 1066 273349 558846 273915
rect 1066 272261 558846 272827
rect 1066 271173 558846 271739
rect 1066 270085 558846 270651
rect 1066 268997 558846 269563
rect 1066 267909 558846 268475
rect 1066 266821 558846 267387
rect 1066 265733 558846 266299
rect 1066 264645 558846 265211
rect 1066 263557 558846 264123
rect 1066 262469 558846 263035
rect 1066 261381 558846 261947
rect 1066 260293 558846 260859
rect 1066 259205 558846 259771
rect 1066 258117 558846 258683
rect 1066 257029 558846 257595
rect 1066 255941 558846 256507
rect 1066 254853 558846 255419
rect 1066 253765 558846 254331
rect 1066 252677 558846 253243
rect 1066 251589 558846 252155
rect 1066 250501 558846 251067
rect 1066 249413 558846 249979
rect 1066 248325 558846 248891
rect 1066 247237 558846 247803
rect 1066 246149 558846 246715
rect 1066 245061 558846 245627
rect 1066 243973 558846 244539
rect 1066 242885 558846 243451
rect 1066 241797 558846 242363
rect 1066 240709 558846 241275
rect 1066 239621 558846 240187
rect 1066 238533 558846 239099
rect 1066 237445 558846 238011
rect 1066 236357 558846 236923
rect 1066 235269 558846 235835
rect 1066 234181 558846 234747
rect 1066 233093 558846 233659
rect 1066 232005 558846 232571
rect 1066 230917 558846 231483
rect 1066 229829 558846 230395
rect 1066 228741 558846 229307
rect 1066 227653 558846 228219
rect 1066 226565 558846 227131
rect 1066 225477 558846 226043
rect 1066 224389 558846 224955
rect 1066 223301 558846 223867
rect 1066 222213 558846 222779
rect 1066 221125 558846 221691
rect 1066 220037 558846 220603
rect 1066 218949 558846 219515
rect 1066 217861 558846 218427
rect 1066 216773 558846 217339
rect 1066 215685 558846 216251
rect 1066 214597 558846 215163
rect 1066 213509 558846 214075
rect 1066 212421 558846 212987
rect 1066 211333 558846 211899
rect 1066 210245 558846 210811
rect 1066 209157 558846 209723
rect 1066 208069 558846 208635
rect 1066 206981 558846 207547
rect 1066 205893 558846 206459
rect 1066 204805 558846 205371
rect 1066 203717 558846 204283
rect 1066 202629 558846 203195
rect 1066 201541 558846 202107
rect 1066 200453 558846 201019
rect 1066 199365 558846 199931
rect 1066 198277 558846 198843
rect 1066 197189 558846 197755
rect 1066 196101 558846 196667
rect 1066 195013 558846 195579
rect 1066 193925 558846 194491
rect 1066 192837 558846 193403
rect 1066 191749 558846 192315
rect 1066 190661 558846 191227
rect 1066 189573 558846 190139
rect 1066 188485 558846 189051
rect 1066 187397 558846 187963
rect 1066 186309 558846 186875
rect 1066 185221 558846 185787
rect 1066 184133 558846 184699
rect 1066 183045 558846 183611
rect 1066 181957 558846 182523
rect 1066 180869 558846 181435
rect 1066 179781 558846 180347
rect 1066 178693 558846 179259
rect 1066 177605 558846 178171
rect 1066 176517 558846 177083
rect 1066 175429 558846 175995
rect 1066 174341 558846 174907
rect 1066 173253 558846 173819
rect 1066 172165 558846 172731
rect 1066 171077 558846 171643
rect 1066 169989 558846 170555
rect 1066 168901 558846 169467
rect 1066 167813 558846 168379
rect 1066 166725 558846 167291
rect 1066 165637 558846 166203
rect 1066 164549 558846 165115
rect 1066 163461 558846 164027
rect 1066 162373 558846 162939
rect 1066 161285 558846 161851
rect 1066 160197 558846 160763
rect 1066 159109 558846 159675
rect 1066 158021 558846 158587
rect 1066 156933 558846 157499
rect 1066 155845 558846 156411
rect 1066 154757 558846 155323
rect 1066 153669 558846 154235
rect 1066 152581 558846 153147
rect 1066 151493 558846 152059
rect 1066 150405 558846 150971
rect 1066 149317 558846 149883
rect 1066 148229 558846 148795
rect 1066 147141 558846 147707
rect 1066 146053 558846 146619
rect 1066 144965 558846 145531
rect 1066 143877 558846 144443
rect 1066 142789 558846 143355
rect 1066 141701 558846 142267
rect 1066 140613 558846 141179
rect 1066 139525 558846 140091
rect 1066 138437 558846 139003
rect 1066 137349 558846 137915
rect 1066 136261 558846 136827
rect 1066 135173 558846 135739
rect 1066 134085 558846 134651
rect 1066 132997 558846 133563
rect 1066 131909 558846 132475
rect 1066 130821 558846 131387
rect 1066 129733 558846 130299
rect 1066 128645 558846 129211
rect 1066 127557 558846 128123
rect 1066 126469 558846 127035
rect 1066 125381 558846 125947
rect 1066 124293 558846 124859
rect 1066 123205 558846 123771
rect 1066 122117 558846 122683
rect 1066 121029 558846 121595
rect 1066 119941 558846 120507
rect 1066 118853 558846 119419
rect 1066 117765 558846 118331
rect 1066 116677 558846 117243
rect 1066 115589 558846 116155
rect 1066 114501 558846 115067
rect 1066 113413 558846 113979
rect 1066 112325 558846 112891
rect 1066 111237 558846 111803
rect 1066 110149 558846 110715
rect 1066 109061 558846 109627
rect 1066 107973 558846 108539
rect 1066 106885 558846 107451
rect 1066 105797 558846 106363
rect 1066 104709 558846 105275
rect 1066 103621 558846 104187
rect 1066 102533 558846 103099
rect 1066 101445 558846 102011
rect 1066 100357 558846 100923
rect 1066 99269 558846 99835
rect 1066 98181 558846 98747
rect 1066 97093 558846 97659
rect 1066 96005 558846 96571
rect 1066 94917 558846 95483
rect 1066 93829 558846 94395
rect 1066 92741 558846 93307
rect 1066 91653 558846 92219
rect 1066 90565 558846 91131
rect 1066 89477 558846 90043
rect 1066 88389 558846 88955
rect 1066 87301 558846 87867
rect 1066 86213 558846 86779
rect 1066 85125 558846 85691
rect 1066 84037 558846 84603
rect 1066 82949 558846 83515
rect 1066 81861 558846 82427
rect 1066 80773 558846 81339
rect 1066 79685 558846 80251
rect 1066 78597 558846 79163
rect 1066 77509 558846 78075
rect 1066 76421 558846 76987
rect 1066 75333 558846 75899
rect 1066 74245 558846 74811
rect 1066 73157 558846 73723
rect 1066 72069 558846 72635
rect 1066 70981 558846 71547
rect 1066 69893 558846 70459
rect 1066 68805 558846 69371
rect 1066 67717 558846 68283
rect 1066 66629 558846 67195
rect 1066 65541 558846 66107
rect 1066 64453 558846 65019
rect 1066 63365 558846 63931
rect 1066 62277 558846 62843
rect 1066 61189 558846 61755
rect 1066 60101 558846 60667
rect 1066 59013 558846 59579
rect 1066 57925 558846 58491
rect 1066 56837 558846 57403
rect 1066 55749 558846 56315
rect 1066 54661 558846 55227
rect 1066 53573 558846 54139
rect 1066 52485 558846 53051
rect 1066 51397 558846 51963
rect 1066 50309 558846 50875
rect 1066 49221 558846 49787
rect 1066 48133 558846 48699
rect 1066 47045 558846 47611
rect 1066 45957 558846 46523
rect 1066 44869 558846 45435
rect 1066 43781 558846 44347
rect 1066 42693 558846 43259
rect 1066 41605 558846 42171
rect 1066 40517 558846 41083
rect 1066 39429 558846 39995
rect 1066 38341 558846 38907
rect 1066 37253 558846 37819
rect 1066 36165 558846 36731
rect 1066 35077 558846 35643
rect 1066 33989 558846 34555
rect 1066 32901 558846 33467
rect 1066 31813 558846 32379
rect 1066 30725 558846 31291
rect 1066 29637 558846 30203
rect 1066 28549 558846 29115
rect 1066 27461 558846 28027
rect 1066 26373 558846 26939
rect 1066 25285 558846 25851
rect 1066 24197 558846 24763
rect 1066 23109 558846 23675
rect 1066 22021 558846 22587
rect 1066 20933 558846 21499
rect 1066 19845 558846 20411
rect 1066 18757 558846 19323
rect 1066 17669 558846 18235
rect 1066 16581 558846 17147
rect 1066 15493 558846 16059
rect 1066 14405 558846 14971
rect 1066 13317 558846 13883
rect 1066 12229 558846 12795
rect 1066 11141 558846 11707
rect 1066 10053 558846 10619
rect 1066 8965 558846 9531
rect 1066 7877 558846 8443
rect 1066 6789 558846 7355
rect 1066 5701 558846 6267
rect 1066 4613 558846 5179
rect 1066 3525 558846 4091
rect 1066 2437 558846 3003
<< obsli1 >>
rect 1104 2159 558808 349809
<< obsm1 >>
rect 1104 76 558808 349840
<< metal2 >>
rect 3146 0 3202 800
rect 8574 0 8630 800
rect 14002 0 14058 800
rect 19430 0 19486 800
rect 24858 0 24914 800
rect 30286 0 30342 800
rect 35714 0 35770 800
rect 41142 0 41198 800
rect 46570 0 46626 800
rect 51998 0 52054 800
rect 57426 0 57482 800
rect 62854 0 62910 800
rect 68282 0 68338 800
rect 73710 0 73766 800
rect 79138 0 79194 800
rect 84566 0 84622 800
rect 89994 0 90050 800
rect 95422 0 95478 800
rect 100850 0 100906 800
rect 106278 0 106334 800
rect 111706 0 111762 800
rect 117134 0 117190 800
rect 122562 0 122618 800
rect 127990 0 128046 800
rect 133418 0 133474 800
rect 138846 0 138902 800
rect 144274 0 144330 800
rect 149702 0 149758 800
rect 155130 0 155186 800
rect 160558 0 160614 800
rect 165986 0 166042 800
rect 171414 0 171470 800
rect 176842 0 176898 800
rect 182270 0 182326 800
rect 187698 0 187754 800
rect 193126 0 193182 800
rect 198554 0 198610 800
rect 203982 0 204038 800
rect 209410 0 209466 800
rect 214838 0 214894 800
rect 220266 0 220322 800
rect 225694 0 225750 800
rect 231122 0 231178 800
rect 236550 0 236606 800
rect 241978 0 242034 800
rect 247406 0 247462 800
rect 252834 0 252890 800
rect 258262 0 258318 800
rect 263690 0 263746 800
rect 269118 0 269174 800
rect 274546 0 274602 800
rect 279974 0 280030 800
rect 285402 0 285458 800
rect 290830 0 290886 800
rect 296258 0 296314 800
rect 301686 0 301742 800
rect 307114 0 307170 800
rect 312542 0 312598 800
rect 317970 0 318026 800
rect 323398 0 323454 800
rect 328826 0 328882 800
rect 334254 0 334310 800
rect 339682 0 339738 800
rect 345110 0 345166 800
rect 350538 0 350594 800
rect 355966 0 356022 800
rect 361394 0 361450 800
rect 366822 0 366878 800
rect 372250 0 372306 800
rect 377678 0 377734 800
rect 383106 0 383162 800
rect 388534 0 388590 800
rect 393962 0 394018 800
rect 399390 0 399446 800
rect 404818 0 404874 800
rect 410246 0 410302 800
rect 415674 0 415730 800
rect 421102 0 421158 800
rect 426530 0 426586 800
rect 431958 0 432014 800
rect 437386 0 437442 800
rect 442814 0 442870 800
rect 448242 0 448298 800
rect 453670 0 453726 800
rect 459098 0 459154 800
rect 464526 0 464582 800
rect 469954 0 470010 800
rect 475382 0 475438 800
rect 480810 0 480866 800
rect 486238 0 486294 800
rect 491666 0 491722 800
rect 497094 0 497150 800
rect 502522 0 502578 800
rect 507950 0 508006 800
rect 513378 0 513434 800
rect 518806 0 518862 800
rect 524234 0 524290 800
rect 529662 0 529718 800
rect 535090 0 535146 800
rect 540518 0 540574 800
rect 545946 0 546002 800
rect 551374 0 551430 800
rect 556802 0 556858 800
<< obsm2 >>
rect 4214 856 557482 349829
rect 4214 70 8518 856
rect 8686 70 13946 856
rect 14114 70 19374 856
rect 19542 70 24802 856
rect 24970 70 30230 856
rect 30398 70 35658 856
rect 35826 70 41086 856
rect 41254 70 46514 856
rect 46682 70 51942 856
rect 52110 70 57370 856
rect 57538 70 62798 856
rect 62966 70 68226 856
rect 68394 70 73654 856
rect 73822 70 79082 856
rect 79250 70 84510 856
rect 84678 70 89938 856
rect 90106 70 95366 856
rect 95534 70 100794 856
rect 100962 70 106222 856
rect 106390 70 111650 856
rect 111818 70 117078 856
rect 117246 70 122506 856
rect 122674 70 127934 856
rect 128102 70 133362 856
rect 133530 70 138790 856
rect 138958 70 144218 856
rect 144386 70 149646 856
rect 149814 70 155074 856
rect 155242 70 160502 856
rect 160670 70 165930 856
rect 166098 70 171358 856
rect 171526 70 176786 856
rect 176954 70 182214 856
rect 182382 70 187642 856
rect 187810 70 193070 856
rect 193238 70 198498 856
rect 198666 70 203926 856
rect 204094 70 209354 856
rect 209522 70 214782 856
rect 214950 70 220210 856
rect 220378 70 225638 856
rect 225806 70 231066 856
rect 231234 70 236494 856
rect 236662 70 241922 856
rect 242090 70 247350 856
rect 247518 70 252778 856
rect 252946 70 258206 856
rect 258374 70 263634 856
rect 263802 70 269062 856
rect 269230 70 274490 856
rect 274658 70 279918 856
rect 280086 70 285346 856
rect 285514 70 290774 856
rect 290942 70 296202 856
rect 296370 70 301630 856
rect 301798 70 307058 856
rect 307226 70 312486 856
rect 312654 70 317914 856
rect 318082 70 323342 856
rect 323510 70 328770 856
rect 328938 70 334198 856
rect 334366 70 339626 856
rect 339794 70 345054 856
rect 345222 70 350482 856
rect 350650 70 355910 856
rect 356078 70 361338 856
rect 361506 70 366766 856
rect 366934 70 372194 856
rect 372362 70 377622 856
rect 377790 70 383050 856
rect 383218 70 388478 856
rect 388646 70 393906 856
rect 394074 70 399334 856
rect 399502 70 404762 856
rect 404930 70 410190 856
rect 410358 70 415618 856
rect 415786 70 421046 856
rect 421214 70 426474 856
rect 426642 70 431902 856
rect 432070 70 437330 856
rect 437498 70 442758 856
rect 442926 70 448186 856
rect 448354 70 453614 856
rect 453782 70 459042 856
rect 459210 70 464470 856
rect 464638 70 469898 856
rect 470066 70 475326 856
rect 475494 70 480754 856
rect 480922 70 486182 856
rect 486350 70 491610 856
rect 491778 70 497038 856
rect 497206 70 502466 856
rect 502634 70 507894 856
rect 508062 70 513322 856
rect 513490 70 518750 856
rect 518918 70 524178 856
rect 524346 70 529606 856
rect 529774 70 535034 856
rect 535202 70 540462 856
rect 540630 70 545890 856
rect 546058 70 551318 856
rect 551486 70 556746 856
rect 556914 70 557482 856
<< obsm3 >>
rect 4210 2143 557486 349825
<< metal4 >>
rect 4208 2128 4528 349840
rect 19568 2128 19888 349840
rect 34928 2128 35248 349840
rect 50288 2128 50608 349840
rect 65648 2128 65968 349840
rect 81008 2128 81328 349840
rect 96368 2128 96688 349840
rect 111728 2128 112048 349840
rect 127088 2128 127408 349840
rect 142448 2128 142768 349840
rect 157808 2128 158128 349840
rect 173168 2128 173488 349840
rect 188528 2128 188848 349840
rect 203888 2128 204208 349840
rect 219248 2128 219568 349840
rect 234608 2128 234928 349840
rect 249968 2128 250288 349840
rect 265328 2128 265648 349840
rect 280688 2128 281008 349840
rect 296048 2128 296368 349840
rect 311408 2128 311728 349840
rect 326768 2128 327088 349840
rect 342128 2128 342448 349840
rect 357488 2128 357808 349840
rect 372848 2128 373168 349840
rect 388208 2128 388528 349840
rect 403568 2128 403888 349840
rect 418928 2128 419248 349840
rect 434288 2128 434608 349840
rect 449648 2128 449968 349840
rect 465008 2128 465328 349840
rect 480368 2128 480688 349840
rect 495728 2128 496048 349840
rect 511088 2128 511408 349840
rect 526448 2128 526768 349840
rect 541808 2128 542128 349840
rect 557168 2128 557488 349840
<< labels >>
rlabel metal2 s 30286 0 30342 800 6 addr_o[0]
port 1 nsew signal output
rlabel metal2 s 203982 0 204038 800 6 addr_o[10]
port 2 nsew signal output
rlabel metal2 s 220266 0 220322 800 6 addr_o[11]
port 3 nsew signal output
rlabel metal2 s 236550 0 236606 800 6 addr_o[12]
port 4 nsew signal output
rlabel metal2 s 252834 0 252890 800 6 addr_o[13]
port 5 nsew signal output
rlabel metal2 s 269118 0 269174 800 6 addr_o[14]
port 6 nsew signal output
rlabel metal2 s 285402 0 285458 800 6 addr_o[15]
port 7 nsew signal output
rlabel metal2 s 301686 0 301742 800 6 addr_o[16]
port 8 nsew signal output
rlabel metal2 s 317970 0 318026 800 6 addr_o[17]
port 9 nsew signal output
rlabel metal2 s 334254 0 334310 800 6 addr_o[18]
port 10 nsew signal output
rlabel metal2 s 350538 0 350594 800 6 addr_o[19]
port 11 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 addr_o[1]
port 12 nsew signal output
rlabel metal2 s 366822 0 366878 800 6 addr_o[20]
port 13 nsew signal output
rlabel metal2 s 383106 0 383162 800 6 addr_o[21]
port 14 nsew signal output
rlabel metal2 s 399390 0 399446 800 6 addr_o[22]
port 15 nsew signal output
rlabel metal2 s 415674 0 415730 800 6 addr_o[23]
port 16 nsew signal output
rlabel metal2 s 431958 0 432014 800 6 addr_o[24]
port 17 nsew signal output
rlabel metal2 s 448242 0 448298 800 6 addr_o[25]
port 18 nsew signal output
rlabel metal2 s 464526 0 464582 800 6 addr_o[26]
port 19 nsew signal output
rlabel metal2 s 480810 0 480866 800 6 addr_o[27]
port 20 nsew signal output
rlabel metal2 s 497094 0 497150 800 6 addr_o[28]
port 21 nsew signal output
rlabel metal2 s 513378 0 513434 800 6 addr_o[29]
port 22 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 addr_o[2]
port 23 nsew signal output
rlabel metal2 s 529662 0 529718 800 6 addr_o[30]
port 24 nsew signal output
rlabel metal2 s 545946 0 546002 800 6 addr_o[31]
port 25 nsew signal output
rlabel metal2 s 89994 0 90050 800 6 addr_o[3]
port 26 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 addr_o[4]
port 27 nsew signal output
rlabel metal2 s 122562 0 122618 800 6 addr_o[5]
port 28 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 addr_o[6]
port 29 nsew signal output
rlabel metal2 s 155130 0 155186 800 6 addr_o[7]
port 30 nsew signal output
rlabel metal2 s 171414 0 171470 800 6 addr_o[8]
port 31 nsew signal output
rlabel metal2 s 187698 0 187754 800 6 addr_o[9]
port 32 nsew signal output
rlabel metal2 s 3146 0 3202 800 6 clk
port 33 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 data_i[0]
port 34 nsew signal input
rlabel metal2 s 209410 0 209466 800 6 data_i[10]
port 35 nsew signal input
rlabel metal2 s 225694 0 225750 800 6 data_i[11]
port 36 nsew signal input
rlabel metal2 s 241978 0 242034 800 6 data_i[12]
port 37 nsew signal input
rlabel metal2 s 258262 0 258318 800 6 data_i[13]
port 38 nsew signal input
rlabel metal2 s 274546 0 274602 800 6 data_i[14]
port 39 nsew signal input
rlabel metal2 s 290830 0 290886 800 6 data_i[15]
port 40 nsew signal input
rlabel metal2 s 307114 0 307170 800 6 data_i[16]
port 41 nsew signal input
rlabel metal2 s 323398 0 323454 800 6 data_i[17]
port 42 nsew signal input
rlabel metal2 s 339682 0 339738 800 6 data_i[18]
port 43 nsew signal input
rlabel metal2 s 355966 0 356022 800 6 data_i[19]
port 44 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 data_i[1]
port 45 nsew signal input
rlabel metal2 s 372250 0 372306 800 6 data_i[20]
port 46 nsew signal input
rlabel metal2 s 388534 0 388590 800 6 data_i[21]
port 47 nsew signal input
rlabel metal2 s 404818 0 404874 800 6 data_i[22]
port 48 nsew signal input
rlabel metal2 s 421102 0 421158 800 6 data_i[23]
port 49 nsew signal input
rlabel metal2 s 437386 0 437442 800 6 data_i[24]
port 50 nsew signal input
rlabel metal2 s 453670 0 453726 800 6 data_i[25]
port 51 nsew signal input
rlabel metal2 s 469954 0 470010 800 6 data_i[26]
port 52 nsew signal input
rlabel metal2 s 486238 0 486294 800 6 data_i[27]
port 53 nsew signal input
rlabel metal2 s 502522 0 502578 800 6 data_i[28]
port 54 nsew signal input
rlabel metal2 s 518806 0 518862 800 6 data_i[29]
port 55 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 data_i[2]
port 56 nsew signal input
rlabel metal2 s 535090 0 535146 800 6 data_i[30]
port 57 nsew signal input
rlabel metal2 s 551374 0 551430 800 6 data_i[31]
port 58 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 data_i[3]
port 59 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 data_i[4]
port 60 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 data_i[5]
port 61 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 data_i[6]
port 62 nsew signal input
rlabel metal2 s 160558 0 160614 800 6 data_i[7]
port 63 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 data_i[8]
port 64 nsew signal input
rlabel metal2 s 193126 0 193182 800 6 data_i[9]
port 65 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 data_o[0]
port 66 nsew signal output
rlabel metal2 s 214838 0 214894 800 6 data_o[10]
port 67 nsew signal output
rlabel metal2 s 231122 0 231178 800 6 data_o[11]
port 68 nsew signal output
rlabel metal2 s 247406 0 247462 800 6 data_o[12]
port 69 nsew signal output
rlabel metal2 s 263690 0 263746 800 6 data_o[13]
port 70 nsew signal output
rlabel metal2 s 279974 0 280030 800 6 data_o[14]
port 71 nsew signal output
rlabel metal2 s 296258 0 296314 800 6 data_o[15]
port 72 nsew signal output
rlabel metal2 s 312542 0 312598 800 6 data_o[16]
port 73 nsew signal output
rlabel metal2 s 328826 0 328882 800 6 data_o[17]
port 74 nsew signal output
rlabel metal2 s 345110 0 345166 800 6 data_o[18]
port 75 nsew signal output
rlabel metal2 s 361394 0 361450 800 6 data_o[19]
port 76 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 data_o[1]
port 77 nsew signal output
rlabel metal2 s 377678 0 377734 800 6 data_o[20]
port 78 nsew signal output
rlabel metal2 s 393962 0 394018 800 6 data_o[21]
port 79 nsew signal output
rlabel metal2 s 410246 0 410302 800 6 data_o[22]
port 80 nsew signal output
rlabel metal2 s 426530 0 426586 800 6 data_o[23]
port 81 nsew signal output
rlabel metal2 s 442814 0 442870 800 6 data_o[24]
port 82 nsew signal output
rlabel metal2 s 459098 0 459154 800 6 data_o[25]
port 83 nsew signal output
rlabel metal2 s 475382 0 475438 800 6 data_o[26]
port 84 nsew signal output
rlabel metal2 s 491666 0 491722 800 6 data_o[27]
port 85 nsew signal output
rlabel metal2 s 507950 0 508006 800 6 data_o[28]
port 86 nsew signal output
rlabel metal2 s 524234 0 524290 800 6 data_o[29]
port 87 nsew signal output
rlabel metal2 s 84566 0 84622 800 6 data_o[2]
port 88 nsew signal output
rlabel metal2 s 540518 0 540574 800 6 data_o[30]
port 89 nsew signal output
rlabel metal2 s 556802 0 556858 800 6 data_o[31]
port 90 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 data_o[3]
port 91 nsew signal output
rlabel metal2 s 117134 0 117190 800 6 data_o[4]
port 92 nsew signal output
rlabel metal2 s 133418 0 133474 800 6 data_o[5]
port 93 nsew signal output
rlabel metal2 s 149702 0 149758 800 6 data_o[6]
port 94 nsew signal output
rlabel metal2 s 165986 0 166042 800 6 data_o[7]
port 95 nsew signal output
rlabel metal2 s 182270 0 182326 800 6 data_o[8]
port 96 nsew signal output
rlabel metal2 s 198554 0 198610 800 6 data_o[9]
port 97 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 done
port 98 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 enable
port 99 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 mem_opdone
port 100 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 mem_operation[0]
port 101 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 mem_operation[1]
port 102 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 reset
port 103 nsew signal input
rlabel metal4 s 4208 2128 4528 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 349840 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 349840 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 349840 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 349840 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 349840 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 349840 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 349840 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 349840 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 349840 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 349840 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 349840 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 349840 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 349840 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 349840 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 349840 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 349840 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 349840 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 349840 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 349840 6 vssd1
port 105 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 50641158
string GDS_FILE /home/leviathan/kicp/openlane/Matrix_Multiplication/runs/23_06_03_14_41/results/signoff/Matrix_Multiplication.magic.gds
string GDS_START 23776
<< end >>

